module main

import wsv

fn main() {
	a := wsv.escape_invalid('allo')
	println(a)
}
